** Profile: "SCHEMATIC1-sim"  [ C:\Users\Georgi\Desktop\P1_2023_434E_Mures_Elena_GSD_N15_OrCad\P1_2023_434E_Mures_Elena_GSD_N15_OrCad\Schematics\15n-pspicefiles\schematic1\sim.sim ] 

** Creating circuit file "sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Cadence/SPB_17.2/tools/pspice/library/New folder/BC856B.lib" 
.LIB "C:/Cadence/SPB_17.2/tools/pspice/library/New folder/BC846B.lib" 
.LIB "C:/Cadence/SPB_17.2/tools/pspice/library/New folder/1N4148.lib" 
.LIB "c:/users/georgi/desktop/smls14bet/smls14bet.lib" 
* From [PSPICE NETLIST] section of C:\Users\Georgi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 0.5ms 0 1u SKIPBP 
.TEMP -20 0 120
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
